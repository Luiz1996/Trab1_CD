CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
290 20 30 60 9
-8 63 1374 736
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
-8 63 1374 736
143654930 0
0
6 Title:
5 Name:
0
0
0
49
13 Logic Switch~
5 555 93 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 E3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 300 89 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 E1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 426 89 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 E2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 800 103 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -17 8 -9
7 CarryIN
-23 -30 26 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 969 100 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 891 100 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
9 Inverter~
13 1054 451 0 2 22
0 8 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U17B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 17 0
1 U
9914 0 0
0
0
14 Logic Display~
6 1463 362 0 1 2
13 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
5 Sa�da
-19 -21 16 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
9 Inverter~
13 619 116 0 2 22
0 12 15
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
3549 0 0
0
0
9 Inverter~
13 358 112 0 2 22
0 19 18
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
7931 0 0
0
0
9 3-In AND~
219 687 147 0 4 22
0 18 16 15 25
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 9 0
1 U
9325 0 0
0
0
9 3-In AND~
219 688 210 0 4 22
0 18 16 12 44
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 9 0
1 U
8903 0 0
0
0
9 3-In AND~
219 690 259 0 4 22
0 18 17 15 22
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 9 0
1 U
3834 0 0
0
0
9 3-In AND~
219 691 310 0 4 22
0 18 17 12 24
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 10 0
1 U
3363 0 0
0
0
9 3-In AND~
219 693 360 0 4 22
0 19 16 15 21
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 10 0
1 U
7668 0 0
0
0
9 3-In AND~
219 695 417 0 4 22
0 19 16 12 43
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U10C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 10 0
1 U
4718 0 0
0
0
9 3-In AND~
219 696 753 0 4 22
0 19 17 15 7
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 11 0
1 U
3874 0 0
0
0
9 3-In AND~
219 702 903 0 4 22
0 19 17 12 10
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U11B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 11 0
1 U
6671 0 0
0
0
9 Inverter~
13 484 112 0 2 22
0 17 16
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
3789 0 0
0
0
8 3-In OR~
219 1408 391 0 4 22
0 3 5 4 20
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U16A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 16 0
1 U
4871 0 0
0
0
14 Logic Display~
6 1464 539 0 1 2
13 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
7 CarryOU
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3750 0 0
0
0
8 2-In OR~
219 1282 614 0 3 22
0 7 10 27
0
0 0 624 90
6 74LS32
-21 -24 21 -16
3 U2B
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8778 0 0
0
0
9 2-In AND~
219 1331 843 0 3 22
0 28 10 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U15D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
538 0 0
0
0
8 3-In OR~
219 1243 834 0 4 22
0 30 29 6 28
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U13C
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 13 0
1 U
6843 0 0
0
0
9 2-In AND~
219 1175 880 0 3 22
0 2 9 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U15C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
3136 0 0
0
0
9 2-In AND~
219 1175 834 0 3 22
0 2 11 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U15B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
5950 0 0
0
0
9 2-In AND~
219 1174 786 0 3 22
0 11 9 30
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U15A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
5670 0 0
0
0
9 2-In AND~
219 1333 703 0 3 22
0 13 7 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
6828 0 0
0
0
9 2-In AND~
219 1331 556 0 3 22
0 31 27 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
6735 0 0
0
0
8 3-In OR~
219 1236 547 0 4 22
0 34 33 32 31
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U13B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 13 0
1 U
8365 0 0
0
0
9 2-In XOR~
219 1180 694 0 3 22
0 35 11 13
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
4132 0 0
0
0
9 2-In XOR~
219 1111 685 0 3 22
0 8 9 35
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
4551 0 0
0
0
9 2-In AND~
219 1168 598 0 3 22
0 8 9 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
3635 0 0
0
0
9 2-In AND~
219 1167 546 0 3 22
0 9 11 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3973 0 0
0
0
9 2-In AND~
219 1167 494 0 3 22
0 8 11 34
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3851 0 0
0
0
8 3-In OR~
219 1234 240 0 4 22
0 41 40 39 42
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U13A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 13 0
1 U
8383 0 0
0
0
8 4-In OR~
219 1317 253 0 5 22
0 42 38 37 36 3
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U12A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0
65 0 0 0 2 1 12 0
1 U
9334 0 0
0
0
9 2-In AND~
219 1165 407 0 3 22
0 45 43 36
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
7471 0 0
0
0
9 2-In AND~
219 1163 351 0 3 22
0 46 21 37
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3334 0 0
0
0
9 2-In AND~
219 1162 301 0 3 22
0 47 24 38
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3559 0 0
0
0
9 2-In AND~
219 1162 249 0 3 22
0 23 22 39
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
984 0 0
0
0
9 2-In AND~
219 1161 201 0 3 22
0 48 44 40
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7557 0 0
0
0
9 2-In AND~
219 1159 138 0 3 22
0 49 25 41
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3146 0 0
0
0
10 2-In XNOR~
219 1047 399 0 3 22
0 8 9 45
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
5687 0 0
0
0
9 2-In XOR~
219 1046 342 0 3 22
0 8 9 46
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7939 0 0
0
0
9 2-In NOR~
219 1042 292 0 3 22
0 8 9 47
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3308 0 0
0
0
10 2-In NAND~
219 1052 240 0 3 22
0 8 9 23
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3408 0 0
0
0
8 2-In OR~
219 1040 191 0 3 22
0 8 9 48
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9773 0 0
0
0
9 2-In AND~
219 1048 129 0 3 22
0 8 9 49
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
691 0 0
0
0
108
1 0 2 0 0 4096 0 25 0 0 7 2
1151 871
1075 871
1 0 2 0 0 0 0 26 0 0 7 2
1151 825
1075 825
5 1 3 0 0 8320 0 37 20 0 0 4
1350 253
1372 253
1372 382
1395 382
3 3 4 0 0 8336 0 23 20 0 0 4
1352 843
1384 843
1384 400
1395 400
3 2 5 0 0 8320 0 28 20 0 0 4
1354 703
1371 703
1371 391
1396 391
3 3 6 0 0 8320 0 24 25 0 0 4
1230 843
1226 843
1226 880
1196 880
2 0 2 0 0 4224 0 7 0 0 0 2
1075 451
1075 988
0 0 7 0 0 4096 0 0 0 0 85 2
907 986
907 753
1 0 8 0 0 4096 0 7 0 0 34 2
1039 451
906 451
1 0 8 0 0 0 0 46 0 0 34 2
1029 283
906 283
2 0 9 0 0 4096 0 44 0 0 30 2
1031 408
991 408
2 0 10 0 0 4096 0 22 0 0 13 2
1294 630
1294 852
2 4 10 0 0 12416 0 23 18 0 0 4
1307 852
1294 852
1294 903
723 903
2 0 9 0 0 4096 0 25 0 0 30 2
1151 889
991 889
2 0 11 0 0 4096 0 26 0 0 36 2
1151 843
820 843
2 0 9 0 0 0 0 27 0 0 30 2
1150 795
991 795
1 0 11 0 0 0 0 27 0 0 36 2
1150 777
820 777
3 0 12 0 0 4096 0 16 0 0 60 4
671 426
588 426
588 427
583 427
2 0 7 0 0 0 0 28 0 0 85 2
1309 712
1276 712
2 0 11 0 0 4096 0 31 0 0 36 2
1164 703
820 703
2 0 9 0 0 0 0 32 0 0 30 2
1095 694
991 694
1 0 8 0 0 4096 0 32 0 0 34 4
1095 676
920 676
920 677
906 677
2 0 9 0 0 0 0 33 0 0 30 2
1144 607
991 607
1 0 8 0 0 4096 0 33 0 0 34 2
1144 589
906 589
2 0 11 0 0 0 0 34 0 0 36 2
1143 555
820 555
1 0 9 0 0 0 0 34 0 0 30 2
1143 537
991 537
2 0 11 0 0 0 0 35 0 0 36 2
1143 503
820 503
1 0 8 0 0 0 0 35 0 0 34 2
1143 485
906 485
1 3 13 0 0 4224 0 28 31 0 0 2
1309 694
1213 694
2 1 9 0 0 4224 0 0 5 0 0 3
991 981
991 100
981 100
0 0 14 0 0 4224 0 0 0 0 0 2
991 100
991 981
1 0 8 0 0 0 0 44 0 0 34 2
1031 390
906 390
1 0 8 0 0 0 0 6 0 0 34 2
903 100
906 100
1 0 8 0 0 8320 0 0 0 33 0 4
903 100
906 100
906 950
907 950
1 0 11 0 0 0 0 4 0 0 36 2
812 103
820 103
1 2 11 0 0 8320 0 0 0 35 0 3
813 103
820 103
820 984
0 3 12 0 0 4096 0 0 18 60 0 2
583 912
678 912
3 0 15 0 0 4096 0 17 0 0 63 2
672 762
622 762
3 0 12 0 0 0 0 14 0 0 60 2
667 319
583 319
3 0 12 0 0 0 0 12 0 0 60 2
664 219
583 219
3 0 15 0 0 0 0 15 0 0 63 2
669 369
622 369
3 0 15 0 0 0 0 13 0 0 63 2
666 268
622 268
3 0 15 0 0 0 0 11 0 0 63 2
663 156
622 156
2 0 16 0 0 4096 0 11 0 0 64 2
663 147
487 147
2 0 16 0 0 4096 0 12 0 0 64 2
664 210
487 210
2 0 17 0 0 4096 0 13 0 0 61 2
666 259
451 259
2 0 17 0 0 4096 0 14 0 0 61 2
667 310
451 310
2 0 16 0 0 4096 0 15 0 0 64 2
669 360
487 360
2 0 16 0 0 0 0 16 0 0 64 4
671 417
502 417
502 416
487 416
2 0 17 0 0 4096 0 17 0 0 61 2
672 753
451 753
2 0 17 0 0 4096 0 18 0 0 61 2
678 903
451 903
1 0 18 0 0 4096 0 11 0 0 65 2
663 138
361 138
1 0 18 0 0 4096 0 12 0 0 65 2
664 201
361 201
1 0 18 0 0 4096 0 13 0 0 65 2
666 250
361 250
1 0 18 0 0 4096 0 14 0 0 65 2
667 301
361 301
1 0 19 0 0 4096 0 15 0 0 62 2
669 351
325 351
1 0 19 0 0 4096 0 16 0 0 62 2
671 408
325 408
1 0 19 0 0 4096 0 17 0 0 62 2
672 744
325 744
1 0 19 0 0 4096 0 18 0 0 62 2
678 894
325 894
1 2 12 0 0 8320 0 0 0 67 0 3
570 92
583 92
583 973
1 2 17 0 0 8320 0 0 0 83 0 3
438 88
451 88
451 969
1 0 19 0 0 8320 0 2 0 0 0 3
312 89
325 89
325 970
2 0 15 0 0 4224 0 9 0 0 0 2
622 134
622 968
2 0 16 0 0 4224 0 19 0 0 0 2
487 130
487 966
2 0 18 0 0 4224 0 10 0 0 0 2
361 130
361 966
4 1 20 0 0 4224 0 20 8 0 0 3
1441 391
1463 391
1463 380
1 1 12 0 0 0 0 1 9 0 0 4
567 93
567 92
622 92
622 98
1 1 19 0 0 0 0 2 10 0 0 4
312 89
312 88
361 88
361 94
2 0 9 0 0 0 0 46 0 0 30 2
1029 301
991 301
1 0 8 0 0 0 0 45 0 0 34 2
1030 333
906 333
2 0 9 0 0 0 0 45 0 0 30 4
1030 351
1010 351
1010 352
991 352
2 4 21 0 0 4224 0 39 15 0 0 2
1139 360
714 360
2 4 22 0 0 12416 0 41 13 0 0 4
1138 258
1109 258
1109 259
711 259
1 3 23 0 0 4224 0 41 47 0 0 2
1138 240
1079 240
2 0 9 0 0 0 0 47 0 0 30 2
1028 249
991 249
1 0 8 0 0 0 0 47 0 0 34 2
1028 231
906 231
2 4 24 0 0 4224 0 40 14 0 0 2
1138 310
712 310
2 0 9 0 0 0 0 49 0 0 30 2
1024 138
991 138
2 0 9 0 0 0 0 48 0 0 30 2
1027 200
991 200
1 0 8 0 0 0 0 48 0 0 34 4
1027 182
929 182
929 181
906 181
1 0 8 0 0 0 0 49 0 0 34 2
1024 120
906 120
2 4 25 0 0 4224 0 43 11 0 0 2
1135 147
708 147
1 1 17 0 0 0 0 3 19 0 0 4
438 89
438 88
487 88
487 94
1 3 26 0 0 8320 0 21 29 0 0 3
1464 557
1464 556
1352 556
4 1 7 0 0 4224 0 17 22 0 0 3
717 753
1276 753
1276 630
2 3 27 0 0 4224 0 29 22 0 0 3
1307 565
1285 565
1285 584
4 1 28 0 0 4224 0 24 23 0 0 2
1276 834
1307 834
2 3 29 0 0 4224 0 24 26 0 0 2
1231 834
1196 834
1 3 30 0 0 4224 0 24 27 0 0 3
1230 825
1230 786
1195 786
4 1 31 0 0 4224 0 30 29 0 0 2
1269 547
1307 547
3 3 32 0 0 8320 0 33 30 0 0 3
1189 598
1223 598
1223 556
2 3 33 0 0 4224 0 30 34 0 0 3
1224 547
1188 547
1188 546
3 1 34 0 0 8320 0 35 30 0 0 3
1188 494
1223 494
1223 538
3 1 35 0 0 4224 0 32 31 0 0 2
1144 685
1164 685
4 3 36 0 0 8320 0 37 38 0 0 4
1300 267
1285 267
1285 407
1186 407
3 3 37 0 0 8320 0 37 39 0 0 4
1300 258
1275 258
1275 351
1184 351
3 2 38 0 0 4224 0 40 37 0 0 4
1183 301
1265 301
1265 249
1300 249
3 3 39 0 0 4224 0 36 41 0 0 2
1221 249
1183 249
2 3 40 0 0 8320 0 36 42 0 0 4
1222 240
1198 240
1198 201
1182 201
1 3 41 0 0 8320 0 36 43 0 0 4
1221 231
1209 231
1209 138
1180 138
4 1 42 0 0 4224 0 36 37 0 0 2
1267 240
1300 240
2 4 43 0 0 8320 0 38 16 0 0 3
1141 416
1141 417
716 417
2 4 44 0 0 4224 0 42 12 0 0 2
1137 210
709 210
3 1 45 0 0 4224 0 44 38 0 0 3
1086 399
1141 399
1141 398
3 1 46 0 0 4224 0 45 39 0 0 2
1079 342
1139 342
3 1 47 0 0 4224 0 46 40 0 0 2
1081 292
1138 292
3 1 48 0 0 4224 0 48 42 0 0 4
1073 191
1118 191
1118 192
1137 192
3 1 49 0 0 4224 0 49 43 0 0 2
1069 129
1135 129
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
858 32 929 51
875 45 938 58
8 ENTRADAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
1003 73 1131 92
1020 86 1140 99
15 FUN��ES L�GICAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
361 22 546 41
377 35 554 48
22          DECODIFICADOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1062 625 1198 644
1079 638 1207 651
16 SOMADOR COMPLETO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
1060 712 1211 731
1076 726 1219 739
18 SUBTRATOR COMPLETO
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
